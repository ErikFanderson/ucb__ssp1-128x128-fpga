parameter NumInstChains = 8;
parameter InstChainLength = 28;
parameter AddressChainLength = 28;
parameter ScanClkDiv = 4;
parameter UARTDataSize = 8;
parameter BaudRate = 256000;
parameter SysClockFrequency = 200000000;

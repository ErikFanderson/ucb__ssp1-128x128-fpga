`default_nettype none
`timescale 1ns/1ps
module ssp1_controller_uart #(
    parameter BaudRate = 9600,
    parameter SystemClockFrequency = 156250000
) (
    input wire i_clk,
    input wire i_rst,
    output wire o_uart_tx,
    input wire i_uart_rx,
    output wire o_uart_rts_n,
    input wire i_uart_cts_n,
    output wire o_mem_reset,
    output wire [7:0] o_mem_leds,
    output wire o_mem_shifter_oe_n,
    output wire o_mem_scan_cg_en,
    input wire [27:0] i_mem_loopback_so_data_0,
    input wire [27:0] i_mem_loopback_so_data_1,
    input wire [27:0] i_mem_loopback_so_data_2,
    input wire [27:0] i_mem_loopback_so_data_3,
    output wire [1:0] o_mem_scan_in_addr_address_0_r0,
    output wire [3:0] o_mem_scan_in_addr_lb_sel_0_r0,
    output wire o_mem_scan_in_addr_enable_0_r0,
    output wire [1:0] o_mem_scan_in_addr_address_0_r1,
    output wire [3:0] o_mem_scan_in_addr_lb_sel_0_r1,
    output wire o_mem_scan_in_addr_enable_0_r1,
    output wire [1:0] o_mem_scan_in_addr_address_0_r2,
    output wire [3:0] o_mem_scan_in_addr_lb_sel_0_r2,
    output wire o_mem_scan_in_addr_enable_0_r2,
    output wire [1:0] o_mem_scan_in_addr_address_0_r3,
    output wire [3:0] o_mem_scan_in_addr_lb_sel_0_r3,
    output wire o_mem_scan_in_addr_enable_0_r3,
    output wire o_mem_scan_in_addr_req_0,
    input wire i_mem_scan_in_addr_ack_0,
    output wire [1:0] o_mem_scan_in_addr_cmd_0,
    output wire [1:0] o_mem_scan_in_addr_address_1_r0,
    output wire [3:0] o_mem_scan_in_addr_lb_sel_1_r0,
    output wire o_mem_scan_in_addr_enable_1_r0,
    output wire [1:0] o_mem_scan_in_addr_address_1_r1,
    output wire [3:0] o_mem_scan_in_addr_lb_sel_1_r1,
    output wire o_mem_scan_in_addr_enable_1_r1,
    output wire [1:0] o_mem_scan_in_addr_address_1_r2,
    output wire [3:0] o_mem_scan_in_addr_lb_sel_1_r2,
    output wire o_mem_scan_in_addr_enable_1_r2,
    output wire [1:0] o_mem_scan_in_addr_address_1_r3,
    output wire [3:0] o_mem_scan_in_addr_lb_sel_1_r3,
    output wire o_mem_scan_in_addr_enable_1_r3,
    output wire o_mem_scan_in_addr_req_1,
    input wire i_mem_scan_in_addr_ack_1,
    output wire [1:0] o_mem_scan_in_addr_cmd_1,
    output wire [1:0] o_mem_scan_in_addr_address_2_r0,
    output wire [3:0] o_mem_scan_in_addr_lb_sel_2_r0,
    output wire o_mem_scan_in_addr_enable_2_r0,
    output wire [1:0] o_mem_scan_in_addr_address_2_r1,
    output wire [3:0] o_mem_scan_in_addr_lb_sel_2_r1,
    output wire o_mem_scan_in_addr_enable_2_r1,
    output wire [1:0] o_mem_scan_in_addr_address_2_r2,
    output wire [3:0] o_mem_scan_in_addr_lb_sel_2_r2,
    output wire o_mem_scan_in_addr_enable_2_r2,
    output wire [1:0] o_mem_scan_in_addr_address_2_r3,
    output wire [3:0] o_mem_scan_in_addr_lb_sel_2_r3,
    output wire o_mem_scan_in_addr_enable_2_r3,
    output wire o_mem_scan_in_addr_req_2,
    input wire i_mem_scan_in_addr_ack_2,
    output wire [1:0] o_mem_scan_in_addr_cmd_2,
    output wire [1:0] o_mem_scan_in_addr_address_3_r0,
    output wire [3:0] o_mem_scan_in_addr_lb_sel_3_r0,
    output wire o_mem_scan_in_addr_enable_3_r0,
    output wire [1:0] o_mem_scan_in_addr_address_3_r1,
    output wire [3:0] o_mem_scan_in_addr_lb_sel_3_r1,
    output wire o_mem_scan_in_addr_enable_3_r1,
    output wire [1:0] o_mem_scan_in_addr_address_3_r2,
    output wire [3:0] o_mem_scan_in_addr_lb_sel_3_r2,
    output wire o_mem_scan_in_addr_enable_3_r2,
    output wire [1:0] o_mem_scan_in_addr_address_3_r3,
    output wire [3:0] o_mem_scan_in_addr_lb_sel_3_r3,
    output wire o_mem_scan_in_addr_enable_3_r3,
    output wire o_mem_scan_in_addr_req_3,
    input wire i_mem_scan_in_addr_ack_3,
    output wire [1:0] o_mem_scan_in_addr_cmd_3,
    output wire [6:0] o_mem_scan_in_inst_0_data_0,
    output wire [6:0] o_mem_scan_in_inst_1_data_0,
    output wire [6:0] o_mem_scan_in_inst_2_data_0,
    output wire [6:0] o_mem_scan_in_inst_3_data_0,
    output wire [6:0] o_mem_scan_in_inst_4_data_0,
    output wire [6:0] o_mem_scan_in_inst_5_data_0,
    output wire [6:0] o_mem_scan_in_inst_6_data_0,
    output wire [6:0] o_mem_scan_in_inst_7_data_0,
    output wire [6:0] o_mem_scan_in_inst_8_data_0,
    output wire [6:0] o_mem_scan_in_inst_9_data_0,
    output wire [6:0] o_mem_scan_in_inst_10_data_0,
    output wire [6:0] o_mem_scan_in_inst_11_data_0,
    output wire [6:0] o_mem_scan_in_inst_12_data_0,
    output wire [6:0] o_mem_scan_in_inst_13_data_0,
    output wire [6:0] o_mem_scan_in_inst_14_data_0,
    output wire [6:0] o_mem_scan_in_inst_15_data_0,
    output wire [6:0] o_mem_scan_in_inst_16_data_0,
    output wire [6:0] o_mem_scan_in_inst_17_data_0,
    output wire [6:0] o_mem_scan_in_inst_18_data_0,
    output wire [6:0] o_mem_scan_in_inst_19_data_0,
    output wire [6:0] o_mem_scan_in_inst_20_data_0,
    output wire [6:0] o_mem_scan_in_inst_21_data_0,
    output wire [6:0] o_mem_scan_in_inst_22_data_0,
    output wire [6:0] o_mem_scan_in_inst_23_data_0,
    output wire [6:0] o_mem_scan_in_inst_24_data_0,
    output wire [6:0] o_mem_scan_in_inst_25_data_0,
    output wire [6:0] o_mem_scan_in_inst_26_data_0,
    output wire [6:0] o_mem_scan_in_inst_27_data_0,
    output wire [6:0] o_mem_scan_in_inst_28_data_0,
    output wire [6:0] o_mem_scan_in_inst_29_data_0,
    output wire [6:0] o_mem_scan_in_inst_30_data_0,
    output wire [6:0] o_mem_scan_in_inst_31_data_0,
    output wire o_mem_scan_in_inst_req_0,
    input wire i_mem_scan_in_inst_ack_0,
    output wire [1:0] o_mem_scan_in_inst_cmd_0,
    output wire [6:0] o_mem_scan_in_inst_0_data_1,
    output wire [6:0] o_mem_scan_in_inst_1_data_1,
    output wire [6:0] o_mem_scan_in_inst_2_data_1,
    output wire [6:0] o_mem_scan_in_inst_3_data_1,
    output wire [6:0] o_mem_scan_in_inst_4_data_1,
    output wire [6:0] o_mem_scan_in_inst_5_data_1,
    output wire [6:0] o_mem_scan_in_inst_6_data_1,
    output wire [6:0] o_mem_scan_in_inst_7_data_1,
    output wire [6:0] o_mem_scan_in_inst_8_data_1,
    output wire [6:0] o_mem_scan_in_inst_9_data_1,
    output wire [6:0] o_mem_scan_in_inst_10_data_1,
    output wire [6:0] o_mem_scan_in_inst_11_data_1,
    output wire [6:0] o_mem_scan_in_inst_12_data_1,
    output wire [6:0] o_mem_scan_in_inst_13_data_1,
    output wire [6:0] o_mem_scan_in_inst_14_data_1,
    output wire [6:0] o_mem_scan_in_inst_15_data_1,
    output wire [6:0] o_mem_scan_in_inst_16_data_1,
    output wire [6:0] o_mem_scan_in_inst_17_data_1,
    output wire [6:0] o_mem_scan_in_inst_18_data_1,
    output wire [6:0] o_mem_scan_in_inst_19_data_1,
    output wire [6:0] o_mem_scan_in_inst_20_data_1,
    output wire [6:0] o_mem_scan_in_inst_21_data_1,
    output wire [6:0] o_mem_scan_in_inst_22_data_1,
    output wire [6:0] o_mem_scan_in_inst_23_data_1,
    output wire [6:0] o_mem_scan_in_inst_24_data_1,
    output wire [6:0] o_mem_scan_in_inst_25_data_1,
    output wire [6:0] o_mem_scan_in_inst_26_data_1,
    output wire [6:0] o_mem_scan_in_inst_27_data_1,
    output wire [6:0] o_mem_scan_in_inst_28_data_1,
    output wire [6:0] o_mem_scan_in_inst_29_data_1,
    output wire [6:0] o_mem_scan_in_inst_30_data_1,
    output wire [6:0] o_mem_scan_in_inst_31_data_1,
    output wire o_mem_scan_in_inst_req_1,
    input wire i_mem_scan_in_inst_ack_1,
    output wire [1:0] o_mem_scan_in_inst_cmd_1,
    output wire [6:0] o_mem_scan_in_inst_0_data_2,
    output wire [6:0] o_mem_scan_in_inst_1_data_2,
    output wire [6:0] o_mem_scan_in_inst_2_data_2,
    output wire [6:0] o_mem_scan_in_inst_3_data_2,
    output wire [6:0] o_mem_scan_in_inst_4_data_2,
    output wire [6:0] o_mem_scan_in_inst_5_data_2,
    output wire [6:0] o_mem_scan_in_inst_6_data_2,
    output wire [6:0] o_mem_scan_in_inst_7_data_2,
    output wire [6:0] o_mem_scan_in_inst_8_data_2,
    output wire [6:0] o_mem_scan_in_inst_9_data_2,
    output wire [6:0] o_mem_scan_in_inst_10_data_2,
    output wire [6:0] o_mem_scan_in_inst_11_data_2,
    output wire [6:0] o_mem_scan_in_inst_12_data_2,
    output wire [6:0] o_mem_scan_in_inst_13_data_2,
    output wire [6:0] o_mem_scan_in_inst_14_data_2,
    output wire [6:0] o_mem_scan_in_inst_15_data_2,
    output wire [6:0] o_mem_scan_in_inst_16_data_2,
    output wire [6:0] o_mem_scan_in_inst_17_data_2,
    output wire [6:0] o_mem_scan_in_inst_18_data_2,
    output wire [6:0] o_mem_scan_in_inst_19_data_2,
    output wire [6:0] o_mem_scan_in_inst_20_data_2,
    output wire [6:0] o_mem_scan_in_inst_21_data_2,
    output wire [6:0] o_mem_scan_in_inst_22_data_2,
    output wire [6:0] o_mem_scan_in_inst_23_data_2,
    output wire [6:0] o_mem_scan_in_inst_24_data_2,
    output wire [6:0] o_mem_scan_in_inst_25_data_2,
    output wire [6:0] o_mem_scan_in_inst_26_data_2,
    output wire [6:0] o_mem_scan_in_inst_27_data_2,
    output wire [6:0] o_mem_scan_in_inst_28_data_2,
    output wire [6:0] o_mem_scan_in_inst_29_data_2,
    output wire [6:0] o_mem_scan_in_inst_30_data_2,
    output wire [6:0] o_mem_scan_in_inst_31_data_2,
    output wire o_mem_scan_in_inst_req_2,
    input wire i_mem_scan_in_inst_ack_2,
    output wire [1:0] o_mem_scan_in_inst_cmd_2,
    output wire [6:0] o_mem_scan_in_inst_0_data_3,
    output wire [6:0] o_mem_scan_in_inst_1_data_3,
    output wire [6:0] o_mem_scan_in_inst_2_data_3,
    output wire [6:0] o_mem_scan_in_inst_3_data_3,
    output wire [6:0] o_mem_scan_in_inst_4_data_3,
    output wire [6:0] o_mem_scan_in_inst_5_data_3,
    output wire [6:0] o_mem_scan_in_inst_6_data_3,
    output wire [6:0] o_mem_scan_in_inst_7_data_3,
    output wire [6:0] o_mem_scan_in_inst_8_data_3,
    output wire [6:0] o_mem_scan_in_inst_9_data_3,
    output wire [6:0] o_mem_scan_in_inst_10_data_3,
    output wire [6:0] o_mem_scan_in_inst_11_data_3,
    output wire [6:0] o_mem_scan_in_inst_12_data_3,
    output wire [6:0] o_mem_scan_in_inst_13_data_3,
    output wire [6:0] o_mem_scan_in_inst_14_data_3,
    output wire [6:0] o_mem_scan_in_inst_15_data_3,
    output wire [6:0] o_mem_scan_in_inst_16_data_3,
    output wire [6:0] o_mem_scan_in_inst_17_data_3,
    output wire [6:0] o_mem_scan_in_inst_18_data_3,
    output wire [6:0] o_mem_scan_in_inst_19_data_3,
    output wire [6:0] o_mem_scan_in_inst_20_data_3,
    output wire [6:0] o_mem_scan_in_inst_21_data_3,
    output wire [6:0] o_mem_scan_in_inst_22_data_3,
    output wire [6:0] o_mem_scan_in_inst_23_data_3,
    output wire [6:0] o_mem_scan_in_inst_24_data_3,
    output wire [6:0] o_mem_scan_in_inst_25_data_3,
    output wire [6:0] o_mem_scan_in_inst_26_data_3,
    output wire [6:0] o_mem_scan_in_inst_27_data_3,
    output wire [6:0] o_mem_scan_in_inst_28_data_3,
    output wire [6:0] o_mem_scan_in_inst_29_data_3,
    output wire [6:0] o_mem_scan_in_inst_30_data_3,
    output wire [6:0] o_mem_scan_in_inst_31_data_3,
    output wire o_mem_scan_in_inst_req_3,
    input wire i_mem_scan_in_inst_ack_3,
    output wire [1:0] o_mem_scan_in_inst_cmd_3,
    output wire o_mem_i2c_req,
    input wire i_mem_i2c_ack,
    output wire [6:0] o_mem_i2c_slave_address,
    output wire [1:0] o_mem_i2c_burst_count_wr,
    output wire [1:0] o_mem_i2c_burst_count_rd,
    output wire [7:0] o_mem_i2c_wdata0,
    output wire [7:0] o_mem_i2c_wdata1,
    output wire [7:0] o_mem_i2c_wdata2,
    output wire [7:0] o_mem_i2c_wdata3,
    output wire o_mem_i2c_rd_wrn,
    input wire i_mem_i2c_nack,
    input wire [7:0] i_mem_i2c_rdata0,
    input wire [7:0] i_mem_i2c_rdata1,
    input wire [7:0] i_mem_i2c_rdata2,
    input wire [7:0] i_mem_i2c_rdata3
);

//--------------------------------------------------------------------------------
// Signals
//--------------------------------------------------------------------------------
wire [7:0] wmem [255:0];
wire [7:0] rmem [255:0];
wire tx_valid;
wire tx_ready;
wire [7:0] tx_data;
wire rx_valid;
wire rx_ready;
wire [7:0] rx_data;
//--------------------------------------------------------------------------------

//--------------------------------------------------------------------------------
// Module instances
//--------------------------------------------------------------------------------
uart #(
    .BaudRate(BaudRate),
    .SystemClockFrequency(SystemClockFrequency),
    .DataSize(8)
) uart_inst (
    .i_clk(i_clk),
    .i_rst(i_rst),
    .i_rx(i_uart_rx),
    .o_tx(o_uart_tx),
    .i_cts_n(i_uart_cts_n),
    .o_rts_n(o_uart_rts_n),
    .o_tx_ready(tx_ready),
    .i_tx_valid(tx_valid),
    .i_tx_data(tx_data),
    .i_rx_ready(rx_ready),
    .o_rx_valid(rx_valid),
    .o_rx_data(rx_data)
);
ssp1_controller_uart_mem_map ssp1_controller_uart_mem_map_inst (
    .ssp1_controller_uart_write_mem(wmem),
    .ssp1_controller_uart_read_mem(rmem),
    .reset(o_mem_reset),
    .leds(o_mem_leds),
    .shifter_oe_n(o_mem_shifter_oe_n),
    .scan_cg_en(o_mem_scan_cg_en),
    .loopback_so_data_0(i_mem_loopback_so_data_0),
    .loopback_so_data_1(i_mem_loopback_so_data_1),
    .loopback_so_data_2(i_mem_loopback_so_data_2),
    .loopback_so_data_3(i_mem_loopback_so_data_3),
    .scan_in_addr_address_0_r0(o_mem_scan_in_addr_address_0_r0),
    .scan_in_addr_lb_sel_0_r0(o_mem_scan_in_addr_lb_sel_0_r0),
    .scan_in_addr_enable_0_r0(o_mem_scan_in_addr_enable_0_r0),
    .scan_in_addr_address_0_r1(o_mem_scan_in_addr_address_0_r1),
    .scan_in_addr_lb_sel_0_r1(o_mem_scan_in_addr_lb_sel_0_r1),
    .scan_in_addr_enable_0_r1(o_mem_scan_in_addr_enable_0_r1),
    .scan_in_addr_address_0_r2(o_mem_scan_in_addr_address_0_r2),
    .scan_in_addr_lb_sel_0_r2(o_mem_scan_in_addr_lb_sel_0_r2),
    .scan_in_addr_enable_0_r2(o_mem_scan_in_addr_enable_0_r2),
    .scan_in_addr_address_0_r3(o_mem_scan_in_addr_address_0_r3),
    .scan_in_addr_lb_sel_0_r3(o_mem_scan_in_addr_lb_sel_0_r3),
    .scan_in_addr_enable_0_r3(o_mem_scan_in_addr_enable_0_r3),
    .scan_in_addr_req_0(o_mem_scan_in_addr_req_0),
    .scan_in_addr_ack_0(i_mem_scan_in_addr_ack_0),
    .scan_in_addr_cmd_0(o_mem_scan_in_addr_cmd_0),
    .scan_in_addr_address_1_r0(o_mem_scan_in_addr_address_1_r0),
    .scan_in_addr_lb_sel_1_r0(o_mem_scan_in_addr_lb_sel_1_r0),
    .scan_in_addr_enable_1_r0(o_mem_scan_in_addr_enable_1_r0),
    .scan_in_addr_address_1_r1(o_mem_scan_in_addr_address_1_r1),
    .scan_in_addr_lb_sel_1_r1(o_mem_scan_in_addr_lb_sel_1_r1),
    .scan_in_addr_enable_1_r1(o_mem_scan_in_addr_enable_1_r1),
    .scan_in_addr_address_1_r2(o_mem_scan_in_addr_address_1_r2),
    .scan_in_addr_lb_sel_1_r2(o_mem_scan_in_addr_lb_sel_1_r2),
    .scan_in_addr_enable_1_r2(o_mem_scan_in_addr_enable_1_r2),
    .scan_in_addr_address_1_r3(o_mem_scan_in_addr_address_1_r3),
    .scan_in_addr_lb_sel_1_r3(o_mem_scan_in_addr_lb_sel_1_r3),
    .scan_in_addr_enable_1_r3(o_mem_scan_in_addr_enable_1_r3),
    .scan_in_addr_req_1(o_mem_scan_in_addr_req_1),
    .scan_in_addr_ack_1(i_mem_scan_in_addr_ack_1),
    .scan_in_addr_cmd_1(o_mem_scan_in_addr_cmd_1),
    .scan_in_addr_address_2_r0(o_mem_scan_in_addr_address_2_r0),
    .scan_in_addr_lb_sel_2_r0(o_mem_scan_in_addr_lb_sel_2_r0),
    .scan_in_addr_enable_2_r0(o_mem_scan_in_addr_enable_2_r0),
    .scan_in_addr_address_2_r1(o_mem_scan_in_addr_address_2_r1),
    .scan_in_addr_lb_sel_2_r1(o_mem_scan_in_addr_lb_sel_2_r1),
    .scan_in_addr_enable_2_r1(o_mem_scan_in_addr_enable_2_r1),
    .scan_in_addr_address_2_r2(o_mem_scan_in_addr_address_2_r2),
    .scan_in_addr_lb_sel_2_r2(o_mem_scan_in_addr_lb_sel_2_r2),
    .scan_in_addr_enable_2_r2(o_mem_scan_in_addr_enable_2_r2),
    .scan_in_addr_address_2_r3(o_mem_scan_in_addr_address_2_r3),
    .scan_in_addr_lb_sel_2_r3(o_mem_scan_in_addr_lb_sel_2_r3),
    .scan_in_addr_enable_2_r3(o_mem_scan_in_addr_enable_2_r3),
    .scan_in_addr_req_2(o_mem_scan_in_addr_req_2),
    .scan_in_addr_ack_2(i_mem_scan_in_addr_ack_2),
    .scan_in_addr_cmd_2(o_mem_scan_in_addr_cmd_2),
    .scan_in_addr_address_3_r0(o_mem_scan_in_addr_address_3_r0),
    .scan_in_addr_lb_sel_3_r0(o_mem_scan_in_addr_lb_sel_3_r0),
    .scan_in_addr_enable_3_r0(o_mem_scan_in_addr_enable_3_r0),
    .scan_in_addr_address_3_r1(o_mem_scan_in_addr_address_3_r1),
    .scan_in_addr_lb_sel_3_r1(o_mem_scan_in_addr_lb_sel_3_r1),
    .scan_in_addr_enable_3_r1(o_mem_scan_in_addr_enable_3_r1),
    .scan_in_addr_address_3_r2(o_mem_scan_in_addr_address_3_r2),
    .scan_in_addr_lb_sel_3_r2(o_mem_scan_in_addr_lb_sel_3_r2),
    .scan_in_addr_enable_3_r2(o_mem_scan_in_addr_enable_3_r2),
    .scan_in_addr_address_3_r3(o_mem_scan_in_addr_address_3_r3),
    .scan_in_addr_lb_sel_3_r3(o_mem_scan_in_addr_lb_sel_3_r3),
    .scan_in_addr_enable_3_r3(o_mem_scan_in_addr_enable_3_r3),
    .scan_in_addr_req_3(o_mem_scan_in_addr_req_3),
    .scan_in_addr_ack_3(i_mem_scan_in_addr_ack_3),
    .scan_in_addr_cmd_3(o_mem_scan_in_addr_cmd_3),
    .scan_in_inst_0_data_0(o_mem_scan_in_inst_0_data_0),
    .scan_in_inst_1_data_0(o_mem_scan_in_inst_1_data_0),
    .scan_in_inst_2_data_0(o_mem_scan_in_inst_2_data_0),
    .scan_in_inst_3_data_0(o_mem_scan_in_inst_3_data_0),
    .scan_in_inst_4_data_0(o_mem_scan_in_inst_4_data_0),
    .scan_in_inst_5_data_0(o_mem_scan_in_inst_5_data_0),
    .scan_in_inst_6_data_0(o_mem_scan_in_inst_6_data_0),
    .scan_in_inst_7_data_0(o_mem_scan_in_inst_7_data_0),
    .scan_in_inst_8_data_0(o_mem_scan_in_inst_8_data_0),
    .scan_in_inst_9_data_0(o_mem_scan_in_inst_9_data_0),
    .scan_in_inst_10_data_0(o_mem_scan_in_inst_10_data_0),
    .scan_in_inst_11_data_0(o_mem_scan_in_inst_11_data_0),
    .scan_in_inst_12_data_0(o_mem_scan_in_inst_12_data_0),
    .scan_in_inst_13_data_0(o_mem_scan_in_inst_13_data_0),
    .scan_in_inst_14_data_0(o_mem_scan_in_inst_14_data_0),
    .scan_in_inst_15_data_0(o_mem_scan_in_inst_15_data_0),
    .scan_in_inst_16_data_0(o_mem_scan_in_inst_16_data_0),
    .scan_in_inst_17_data_0(o_mem_scan_in_inst_17_data_0),
    .scan_in_inst_18_data_0(o_mem_scan_in_inst_18_data_0),
    .scan_in_inst_19_data_0(o_mem_scan_in_inst_19_data_0),
    .scan_in_inst_20_data_0(o_mem_scan_in_inst_20_data_0),
    .scan_in_inst_21_data_0(o_mem_scan_in_inst_21_data_0),
    .scan_in_inst_22_data_0(o_mem_scan_in_inst_22_data_0),
    .scan_in_inst_23_data_0(o_mem_scan_in_inst_23_data_0),
    .scan_in_inst_24_data_0(o_mem_scan_in_inst_24_data_0),
    .scan_in_inst_25_data_0(o_mem_scan_in_inst_25_data_0),
    .scan_in_inst_26_data_0(o_mem_scan_in_inst_26_data_0),
    .scan_in_inst_27_data_0(o_mem_scan_in_inst_27_data_0),
    .scan_in_inst_28_data_0(o_mem_scan_in_inst_28_data_0),
    .scan_in_inst_29_data_0(o_mem_scan_in_inst_29_data_0),
    .scan_in_inst_30_data_0(o_mem_scan_in_inst_30_data_0),
    .scan_in_inst_31_data_0(o_mem_scan_in_inst_31_data_0),
    .scan_in_inst_req_0(o_mem_scan_in_inst_req_0),
    .scan_in_inst_ack_0(i_mem_scan_in_inst_ack_0),
    .scan_in_inst_cmd_0(o_mem_scan_in_inst_cmd_0),
    .scan_in_inst_0_data_1(o_mem_scan_in_inst_0_data_1),
    .scan_in_inst_1_data_1(o_mem_scan_in_inst_1_data_1),
    .scan_in_inst_2_data_1(o_mem_scan_in_inst_2_data_1),
    .scan_in_inst_3_data_1(o_mem_scan_in_inst_3_data_1),
    .scan_in_inst_4_data_1(o_mem_scan_in_inst_4_data_1),
    .scan_in_inst_5_data_1(o_mem_scan_in_inst_5_data_1),
    .scan_in_inst_6_data_1(o_mem_scan_in_inst_6_data_1),
    .scan_in_inst_7_data_1(o_mem_scan_in_inst_7_data_1),
    .scan_in_inst_8_data_1(o_mem_scan_in_inst_8_data_1),
    .scan_in_inst_9_data_1(o_mem_scan_in_inst_9_data_1),
    .scan_in_inst_10_data_1(o_mem_scan_in_inst_10_data_1),
    .scan_in_inst_11_data_1(o_mem_scan_in_inst_11_data_1),
    .scan_in_inst_12_data_1(o_mem_scan_in_inst_12_data_1),
    .scan_in_inst_13_data_1(o_mem_scan_in_inst_13_data_1),
    .scan_in_inst_14_data_1(o_mem_scan_in_inst_14_data_1),
    .scan_in_inst_15_data_1(o_mem_scan_in_inst_15_data_1),
    .scan_in_inst_16_data_1(o_mem_scan_in_inst_16_data_1),
    .scan_in_inst_17_data_1(o_mem_scan_in_inst_17_data_1),
    .scan_in_inst_18_data_1(o_mem_scan_in_inst_18_data_1),
    .scan_in_inst_19_data_1(o_mem_scan_in_inst_19_data_1),
    .scan_in_inst_20_data_1(o_mem_scan_in_inst_20_data_1),
    .scan_in_inst_21_data_1(o_mem_scan_in_inst_21_data_1),
    .scan_in_inst_22_data_1(o_mem_scan_in_inst_22_data_1),
    .scan_in_inst_23_data_1(o_mem_scan_in_inst_23_data_1),
    .scan_in_inst_24_data_1(o_mem_scan_in_inst_24_data_1),
    .scan_in_inst_25_data_1(o_mem_scan_in_inst_25_data_1),
    .scan_in_inst_26_data_1(o_mem_scan_in_inst_26_data_1),
    .scan_in_inst_27_data_1(o_mem_scan_in_inst_27_data_1),
    .scan_in_inst_28_data_1(o_mem_scan_in_inst_28_data_1),
    .scan_in_inst_29_data_1(o_mem_scan_in_inst_29_data_1),
    .scan_in_inst_30_data_1(o_mem_scan_in_inst_30_data_1),
    .scan_in_inst_31_data_1(o_mem_scan_in_inst_31_data_1),
    .scan_in_inst_req_1(o_mem_scan_in_inst_req_1),
    .scan_in_inst_ack_1(i_mem_scan_in_inst_ack_1),
    .scan_in_inst_cmd_1(o_mem_scan_in_inst_cmd_1),
    .scan_in_inst_0_data_2(o_mem_scan_in_inst_0_data_2),
    .scan_in_inst_1_data_2(o_mem_scan_in_inst_1_data_2),
    .scan_in_inst_2_data_2(o_mem_scan_in_inst_2_data_2),
    .scan_in_inst_3_data_2(o_mem_scan_in_inst_3_data_2),
    .scan_in_inst_4_data_2(o_mem_scan_in_inst_4_data_2),
    .scan_in_inst_5_data_2(o_mem_scan_in_inst_5_data_2),
    .scan_in_inst_6_data_2(o_mem_scan_in_inst_6_data_2),
    .scan_in_inst_7_data_2(o_mem_scan_in_inst_7_data_2),
    .scan_in_inst_8_data_2(o_mem_scan_in_inst_8_data_2),
    .scan_in_inst_9_data_2(o_mem_scan_in_inst_9_data_2),
    .scan_in_inst_10_data_2(o_mem_scan_in_inst_10_data_2),
    .scan_in_inst_11_data_2(o_mem_scan_in_inst_11_data_2),
    .scan_in_inst_12_data_2(o_mem_scan_in_inst_12_data_2),
    .scan_in_inst_13_data_2(o_mem_scan_in_inst_13_data_2),
    .scan_in_inst_14_data_2(o_mem_scan_in_inst_14_data_2),
    .scan_in_inst_15_data_2(o_mem_scan_in_inst_15_data_2),
    .scan_in_inst_16_data_2(o_mem_scan_in_inst_16_data_2),
    .scan_in_inst_17_data_2(o_mem_scan_in_inst_17_data_2),
    .scan_in_inst_18_data_2(o_mem_scan_in_inst_18_data_2),
    .scan_in_inst_19_data_2(o_mem_scan_in_inst_19_data_2),
    .scan_in_inst_20_data_2(o_mem_scan_in_inst_20_data_2),
    .scan_in_inst_21_data_2(o_mem_scan_in_inst_21_data_2),
    .scan_in_inst_22_data_2(o_mem_scan_in_inst_22_data_2),
    .scan_in_inst_23_data_2(o_mem_scan_in_inst_23_data_2),
    .scan_in_inst_24_data_2(o_mem_scan_in_inst_24_data_2),
    .scan_in_inst_25_data_2(o_mem_scan_in_inst_25_data_2),
    .scan_in_inst_26_data_2(o_mem_scan_in_inst_26_data_2),
    .scan_in_inst_27_data_2(o_mem_scan_in_inst_27_data_2),
    .scan_in_inst_28_data_2(o_mem_scan_in_inst_28_data_2),
    .scan_in_inst_29_data_2(o_mem_scan_in_inst_29_data_2),
    .scan_in_inst_30_data_2(o_mem_scan_in_inst_30_data_2),
    .scan_in_inst_31_data_2(o_mem_scan_in_inst_31_data_2),
    .scan_in_inst_req_2(o_mem_scan_in_inst_req_2),
    .scan_in_inst_ack_2(i_mem_scan_in_inst_ack_2),
    .scan_in_inst_cmd_2(o_mem_scan_in_inst_cmd_2),
    .scan_in_inst_0_data_3(o_mem_scan_in_inst_0_data_3),
    .scan_in_inst_1_data_3(o_mem_scan_in_inst_1_data_3),
    .scan_in_inst_2_data_3(o_mem_scan_in_inst_2_data_3),
    .scan_in_inst_3_data_3(o_mem_scan_in_inst_3_data_3),
    .scan_in_inst_4_data_3(o_mem_scan_in_inst_4_data_3),
    .scan_in_inst_5_data_3(o_mem_scan_in_inst_5_data_3),
    .scan_in_inst_6_data_3(o_mem_scan_in_inst_6_data_3),
    .scan_in_inst_7_data_3(o_mem_scan_in_inst_7_data_3),
    .scan_in_inst_8_data_3(o_mem_scan_in_inst_8_data_3),
    .scan_in_inst_9_data_3(o_mem_scan_in_inst_9_data_3),
    .scan_in_inst_10_data_3(o_mem_scan_in_inst_10_data_3),
    .scan_in_inst_11_data_3(o_mem_scan_in_inst_11_data_3),
    .scan_in_inst_12_data_3(o_mem_scan_in_inst_12_data_3),
    .scan_in_inst_13_data_3(o_mem_scan_in_inst_13_data_3),
    .scan_in_inst_14_data_3(o_mem_scan_in_inst_14_data_3),
    .scan_in_inst_15_data_3(o_mem_scan_in_inst_15_data_3),
    .scan_in_inst_16_data_3(o_mem_scan_in_inst_16_data_3),
    .scan_in_inst_17_data_3(o_mem_scan_in_inst_17_data_3),
    .scan_in_inst_18_data_3(o_mem_scan_in_inst_18_data_3),
    .scan_in_inst_19_data_3(o_mem_scan_in_inst_19_data_3),
    .scan_in_inst_20_data_3(o_mem_scan_in_inst_20_data_3),
    .scan_in_inst_21_data_3(o_mem_scan_in_inst_21_data_3),
    .scan_in_inst_22_data_3(o_mem_scan_in_inst_22_data_3),
    .scan_in_inst_23_data_3(o_mem_scan_in_inst_23_data_3),
    .scan_in_inst_24_data_3(o_mem_scan_in_inst_24_data_3),
    .scan_in_inst_25_data_3(o_mem_scan_in_inst_25_data_3),
    .scan_in_inst_26_data_3(o_mem_scan_in_inst_26_data_3),
    .scan_in_inst_27_data_3(o_mem_scan_in_inst_27_data_3),
    .scan_in_inst_28_data_3(o_mem_scan_in_inst_28_data_3),
    .scan_in_inst_29_data_3(o_mem_scan_in_inst_29_data_3),
    .scan_in_inst_30_data_3(o_mem_scan_in_inst_30_data_3),
    .scan_in_inst_31_data_3(o_mem_scan_in_inst_31_data_3),
    .scan_in_inst_req_3(o_mem_scan_in_inst_req_3),
    .scan_in_inst_ack_3(i_mem_scan_in_inst_ack_3),
    .scan_in_inst_cmd_3(o_mem_scan_in_inst_cmd_3),
    .i2c_req(o_mem_i2c_req),
    .i2c_ack(i_mem_i2c_ack),
    .i2c_slave_address(o_mem_i2c_slave_address),
    .i2c_burst_count_wr(o_mem_i2c_burst_count_wr),
    .i2c_burst_count_rd(o_mem_i2c_burst_count_rd),
    .i2c_wdata0(o_mem_i2c_wdata0),
    .i2c_wdata1(o_mem_i2c_wdata1),
    .i2c_wdata2(o_mem_i2c_wdata2),
    .i2c_wdata3(o_mem_i2c_wdata3),
    .i2c_rd_wrn(o_mem_i2c_rd_wrn),
    .i2c_nack(i_mem_i2c_nack),
    .i2c_rdata0(i_mem_i2c_rdata0),
    .i2c_rdata1(i_mem_i2c_rdata1),
    .i2c_rdata2(i_mem_i2c_rdata2),
    .i2c_rdata3(i_mem_i2c_rdata3)
);
uart_mem_access #(
    .DataSize(8),
    .AddressSize(8)
) uart_mem_access_inst (
    .i_clk(i_clk),
    .i_rst(i_rst),
    .i_rx_data(rx_data),
    .i_rx_valid(rx_valid),
    .o_rx_ready(rx_ready),
    .o_tx_data(tx_data),
    .o_tx_valid(tx_valid),
    .i_tx_ready(tx_ready),
    .o_wmem(wmem),
    .i_rmem(rmem)
);
//--------------------------------------------------------------------------------

//--------------------------------------------------------------------------------
// Task declarations
//--------------------------------------------------------------------------------
//--------------------------------------------------------------------------------

//--------------------------------------------------------------------------------
// Initial statements
//--------------------------------------------------------------------------------
//--------------------------------------------------------------------------------

//--------------------------------------------------------------------------------
// Internals of module
//--------------------------------------------------------------------------------
//--------------------------------------------------------------------------------

endmodule
`default_nettype wire

parameter NumInstChains = 8;
parameter InstChainLength = 28;
parameter AddressChainLength = 28;
parameter ScanClkDiv = 128;
parameter UARTDataSize = 8;
parameter BaudRate = 64000;
parameter SysClockFrequency = 156250000;
parameter MaxUserFrequency = 156250000;

//==============================================================================
// Author: Erik Anderson 
// Email: efa@eecs.berkeley.edu
// Description: Top level testbench for "ssp1_controller"
// Naming conventions:
//    signals => snake_case
//    Parameters (aliasing signal values) => SNAKE_CASE with all caps
//    Parameters (not aliasing signal values) => CamelCase 
//==============================================================================

module top;

// Data input interface
wire o_scan_clk_p;
wire o_scan_clk_n;
wire [3:0] o_scan_reset;
wire [3:0] o_scan_update;
wire [3:0] o_scan_en_inst;
wire [3:0] [7:0] o_scan_in_inst;
    
// Data output interface (for debug)
wire [3:0] i_scan_clk_p;
wire [3:0] i_scan_clk_n;
wire [3:0] i_scan_reset;
wire [3:0] i_scan_update;
wire [3:0] i_scan_en_inst;
wire [3:0] [7:0] i_scan_in_inst;

// Address scan in/out and enable signals
wire [3:0] o_scan_in_address;
wire [3:0] i_scan_out_address;
wire [3:0] o_scan_en_address;
wire [3:0] i_scan_en_address;

// Misc signals - loopback debug and level shifter output enable
wire [3:0] o_scan_in_loopback;
wire [3:0] i_scan_out_loopback;

// UART signals
wire uart_tx, uart_rx;
wire uart_cts_n, uart_rts_n;

wire [3:0] [31:0] [31:0] mems_output;
//-----------------------------------------------------------------------------
// Instances
//-----------------------------------------------------------------------------
// Instantiate Bus Functional Model (BFM) interface
ssp1_controller_bfm bfm();
 
// Instantiate Device Under Test (DUT) 
ssp1_controller #(
    .NumInstChains(bfm.NumInstChains),
    .InstChainLength(bfm.InstChainLength),
    .AddressChainLength(bfm.AddressChainLength),
    .ScanClkDiv(bfm.ScanClkDiv), 
    .UARTDataSize(bfm.UARTDataSize),
    .BaudRate(bfm.BaudRate),
    .SysClockFrequency(bfm.SysClockFrequency)
) dut (
    .i_sys_clk(bfm.i_sys_clk),
    .i_user_clk(bfm.i_user_clk),
    .i_rst(bfm.i_rst),
    .o_shifter_oe_n(bfm.o_shifter_oe_n),
    .o_led(bfm.o_led),

    .o_uart_tx(uart_rx),
    .i_uart_rx(uart_tx),
    .o_uart_rts_n(uart_cts_n),
    .i_uart_cts_n(uart_rts_n),

    .i_sda(bfm.i_sda),
    .i_scl(bfm.i_scl),
    .o_sda_oe_n(bfm.o_sda_oe_n),
    .o_scl_oe_n(bfm.o_scl_oe_n),

    .o_scan_clk_p(o_scan_clk_p),
    .o_scan_clk_n(o_scan_clk_n),
    .o_scan_reset(o_scan_reset),
    .o_scan_update(o_scan_update),
    .o_scan_en_inst(o_scan_en_inst),
    .o_scan_in_inst(o_scan_in_inst),
    .o_scan_in_address(o_scan_in_address),
    .o_scan_en_address(o_scan_en_address),
    .i_scan_out_loopback(i_scan_out_loopback)
);

// Instantiate UART that will emulate PC UART
uart #(
    .BaudRate(bfm.BaudRate),
    .SystemClockFrequency(bfm.SysClockFrequency),
    .DataSize(bfm.UARTDataSize)
) uart_inst (
    .i_clk(bfm.i_sys_clk),
    .i_rst(bfm.i_rst),
    
    .i_rx(uart_rx),
    .o_tx(uart_tx),
    .i_cts_n(uart_cts_n),
    .o_rts_n(uart_rts_n),
    
    .o_tx_ready(bfm.tx_ready),
    .i_tx_valid(bfm.tx_valid),
    .i_tx_data(bfm.tx_data),
    .i_rx_ready(bfm.rx_ready),
    .o_rx_valid(bfm.rx_valid),
    .o_rx_data(bfm.rx_data)
);

// Instantiate chip model (leave mems outputs disconnected)
genvar i;
generate for (i = 0; i < 4; i++) begin
    MemsSwitchController chip (
        .io_scanClkPIn(o_scan_clk_p),
        .io_scanClkPOut(i_scan_clk_p[i]),
        .io_scanClkNIn(o_scan_clk_n),
        .io_scanClkNOut(i_scan_clk_n[i]),
        .io_scanUpdateIn(o_scan_update[i]),
        .io_scanUpdateOut(i_scan_update[i]),
        .io_scanResetIn(o_scan_reset[i]),
        .io_scanResetOut(i_scan_reset[i]),
        .io_scanEnInstIn(o_scan_en_inst[i]),
        .io_scanEnInstOut(i_scan_en_inst[i]),
        .io_scanInAddress(o_scan_in_address[i]),
        .io_scanOutAddress(i_scan_out_address[i]),
        .io_scanEnAddressIn(o_scan_en_address[i]),
        .io_scanEnAddressOut(i_scan_en_address[i]),
        .io_scanOutLoopback(i_scan_out_loopback[i]),
        .io_scanInLoopback(o_scan_in_loopback[i]),
        .io_scanInInstIn_0(o_scan_in_inst[i][0]),
        .io_scanInInstOut_0(i_scan_in_inst[i][0]),
        .io_scanInInstIn_1(o_scan_in_inst[i][1]),
        .io_scanInInstOut_1(i_scan_in_inst[i][1]),
        .io_scanInInstIn_2(o_scan_in_inst[i][2]),
        .io_scanInInstOut_2(i_scan_in_inst[i][2]),
        .io_scanInInstIn_3(o_scan_in_inst[i][3]),
        .io_scanInInstOut_3(i_scan_in_inst[i][3]),
        .io_scanInInstIn_4(o_scan_in_inst[i][4]),
        .io_scanInInstOut_4(i_scan_in_inst[i][4]),
        .io_scanInInstIn_5(o_scan_in_inst[i][5]),
        .io_scanInInstOut_5(i_scan_in_inst[i][5]),
        .io_scanInInstIn_6(o_scan_in_inst[i][6]),
        .io_scanInInstOut_6(i_scan_in_inst[i][6]),
        .io_scanInInstIn_7(o_scan_in_inst[i][7]),
        .io_scanInInstOut_7(i_scan_in_inst[i][7]),
        .io_output_0_0(mems_output[i][0][0]),
        .io_output_0_1(mems_output[i][0][1]),
        .io_output_0_2(mems_output[i][0][2]),
        .io_output_0_3(mems_output[i][0][3]),
        .io_output_0_4(mems_output[i][0][4]),
        .io_output_0_5(mems_output[i][0][5]),
        .io_output_0_6(mems_output[i][0][6]),
        .io_output_0_7(mems_output[i][0][7]),
        .io_output_0_8(mems_output[i][0][8]),
        .io_output_0_9(mems_output[i][0][9]),
        .io_output_0_10(mems_output[i][0][10]),
        .io_output_0_11(mems_output[i][0][11]),
        .io_output_0_12(mems_output[i][0][12]),
        .io_output_0_13(mems_output[i][0][13]),
        .io_output_0_14(mems_output[i][0][14]),
        .io_output_0_15(mems_output[i][0][15]),
        .io_output_0_16(mems_output[i][0][16]),
        .io_output_0_17(mems_output[i][0][17]),
        .io_output_0_18(mems_output[i][0][18]),
        .io_output_0_19(mems_output[i][0][19]),
        .io_output_0_20(mems_output[i][0][20]),
        .io_output_0_21(mems_output[i][0][21]),
        .io_output_0_22(mems_output[i][0][22]),
        .io_output_0_23(mems_output[i][0][23]),
        .io_output_0_24(mems_output[i][0][24]),
        .io_output_0_25(mems_output[i][0][25]),
        .io_output_0_26(mems_output[i][0][26]),
        .io_output_0_27(mems_output[i][0][27]),
        .io_output_0_28(mems_output[i][0][28]),
        .io_output_0_29(mems_output[i][0][29]),
        .io_output_0_30(mems_output[i][0][30]),
        .io_output_0_31(mems_output[i][0][31]),
        .io_output_1_0(mems_output[i][1][0]),
        .io_output_1_1(mems_output[i][1][1]),
        .io_output_1_2(mems_output[i][1][2]),
        .io_output_1_3(mems_output[i][1][3]),
        .io_output_1_4(mems_output[i][1][4]),
        .io_output_1_5(mems_output[i][1][5]),
        .io_output_1_6(mems_output[i][1][6]),
        .io_output_1_7(mems_output[i][1][7]),
        .io_output_1_8(mems_output[i][1][8]),
        .io_output_1_9(mems_output[i][1][9]),
        .io_output_1_10(mems_output[i][1][10]),
        .io_output_1_11(mems_output[i][1][11]),
        .io_output_1_12(mems_output[i][1][12]),
        .io_output_1_13(mems_output[i][1][13]),
        .io_output_1_14(mems_output[i][1][14]),
        .io_output_1_15(mems_output[i][1][15]),
        .io_output_1_16(mems_output[i][1][16]),
        .io_output_1_17(mems_output[i][1][17]),
        .io_output_1_18(mems_output[i][1][18]),
        .io_output_1_19(mems_output[i][1][19]),
        .io_output_1_20(mems_output[i][1][20]),
        .io_output_1_21(mems_output[i][1][21]),
        .io_output_1_22(mems_output[i][1][22]),
        .io_output_1_23(mems_output[i][1][23]),
        .io_output_1_24(mems_output[i][1][24]),
        .io_output_1_25(mems_output[i][1][25]),
        .io_output_1_26(mems_output[i][1][26]),
        .io_output_1_27(mems_output[i][1][27]),
        .io_output_1_28(mems_output[i][1][28]),
        .io_output_1_29(mems_output[i][1][29]),
        .io_output_1_30(mems_output[i][1][30]),
        .io_output_1_31(mems_output[i][1][31]),
        .io_output_2_0(mems_output[i][2][0]),
        .io_output_2_1(mems_output[i][2][1]),
        .io_output_2_2(mems_output[i][2][2]),
        .io_output_2_3(mems_output[i][2][3]),
        .io_output_2_4(mems_output[i][2][4]),
        .io_output_2_5(mems_output[i][2][5]),
        .io_output_2_6(mems_output[i][2][6]),
        .io_output_2_7(mems_output[i][2][7]),
        .io_output_2_8(mems_output[i][2][8]),
        .io_output_2_9(mems_output[i][2][9]),
        .io_output_2_10(mems_output[i][2][10]),
        .io_output_2_11(mems_output[i][2][11]),
        .io_output_2_12(mems_output[i][2][12]),
        .io_output_2_13(mems_output[i][2][13]),
        .io_output_2_14(mems_output[i][2][14]),
        .io_output_2_15(mems_output[i][2][15]),
        .io_output_2_16(mems_output[i][2][16]),
        .io_output_2_17(mems_output[i][2][17]),
        .io_output_2_18(mems_output[i][2][18]),
        .io_output_2_19(mems_output[i][2][19]),
        .io_output_2_20(mems_output[i][2][20]),
        .io_output_2_21(mems_output[i][2][21]),
        .io_output_2_22(mems_output[i][2][22]),
        .io_output_2_23(mems_output[i][2][23]),
        .io_output_2_24(mems_output[i][2][24]),
        .io_output_2_25(mems_output[i][2][25]),
        .io_output_2_26(mems_output[i][2][26]),
        .io_output_2_27(mems_output[i][2][27]),
        .io_output_2_28(mems_output[i][2][28]),
        .io_output_2_29(mems_output[i][2][29]),
        .io_output_2_30(mems_output[i][2][30]),
        .io_output_2_31(mems_output[i][2][31]),
        .io_output_3_0(mems_output[i][3][0]),
        .io_output_3_1(mems_output[i][3][1]),
        .io_output_3_2(mems_output[i][3][2]),
        .io_output_3_3(mems_output[i][3][3]),
        .io_output_3_4(mems_output[i][3][4]),
        .io_output_3_5(mems_output[i][3][5]),
        .io_output_3_6(mems_output[i][3][6]),
        .io_output_3_7(mems_output[i][3][7]),
        .io_output_3_8(mems_output[i][3][8]),
        .io_output_3_9(mems_output[i][3][9]),
        .io_output_3_10(mems_output[i][3][10]),
        .io_output_3_11(mems_output[i][3][11]),
        .io_output_3_12(mems_output[i][3][12]),
        .io_output_3_13(mems_output[i][3][13]),
        .io_output_3_14(mems_output[i][3][14]),
        .io_output_3_15(mems_output[i][3][15]),
        .io_output_3_16(mems_output[i][3][16]),
        .io_output_3_17(mems_output[i][3][17]),
        .io_output_3_18(mems_output[i][3][18]),
        .io_output_3_19(mems_output[i][3][19]),
        .io_output_3_20(mems_output[i][3][20]),
        .io_output_3_21(mems_output[i][3][21]),
        .io_output_3_22(mems_output[i][3][22]),
        .io_output_3_23(mems_output[i][3][23]),
        .io_output_3_24(mems_output[i][3][24]),
        .io_output_3_25(mems_output[i][3][25]),
        .io_output_3_26(mems_output[i][3][26]),
        .io_output_3_27(mems_output[i][3][27]),
        .io_output_3_28(mems_output[i][3][28]),
        .io_output_3_29(mems_output[i][3][29]),
        .io_output_3_30(mems_output[i][3][30]),
        .io_output_3_31(mems_output[i][3][31]),
        .io_output_4_0(mems_output[i][4][0]),
        .io_output_4_1(mems_output[i][4][1]),
        .io_output_4_2(mems_output[i][4][2]),
        .io_output_4_3(mems_output[i][4][3]),
        .io_output_4_4(mems_output[i][4][4]),
        .io_output_4_5(mems_output[i][4][5]),
        .io_output_4_6(mems_output[i][4][6]),
        .io_output_4_7(mems_output[i][4][7]),
        .io_output_4_8(mems_output[i][4][8]),
        .io_output_4_9(mems_output[i][4][9]),
        .io_output_4_10(mems_output[i][4][10]),
        .io_output_4_11(mems_output[i][4][11]),
        .io_output_4_12(mems_output[i][4][12]),
        .io_output_4_13(mems_output[i][4][13]),
        .io_output_4_14(mems_output[i][4][14]),
        .io_output_4_15(mems_output[i][4][15]),
        .io_output_4_16(mems_output[i][4][16]),
        .io_output_4_17(mems_output[i][4][17]),
        .io_output_4_18(mems_output[i][4][18]),
        .io_output_4_19(mems_output[i][4][19]),
        .io_output_4_20(mems_output[i][4][20]),
        .io_output_4_21(mems_output[i][4][21]),
        .io_output_4_22(mems_output[i][4][22]),
        .io_output_4_23(mems_output[i][4][23]),
        .io_output_4_24(mems_output[i][4][24]),
        .io_output_4_25(mems_output[i][4][25]),
        .io_output_4_26(mems_output[i][4][26]),
        .io_output_4_27(mems_output[i][4][27]),
        .io_output_4_28(mems_output[i][4][28]),
        .io_output_4_29(mems_output[i][4][29]),
        .io_output_4_30(mems_output[i][4][30]),
        .io_output_4_31(mems_output[i][4][31]),
        .io_output_5_0(mems_output[i][5][0]),
        .io_output_5_1(mems_output[i][5][1]),
        .io_output_5_2(mems_output[i][5][2]),
        .io_output_5_3(mems_output[i][5][3]),
        .io_output_5_4(mems_output[i][5][4]),
        .io_output_5_5(mems_output[i][5][5]),
        .io_output_5_6(mems_output[i][5][6]),
        .io_output_5_7(mems_output[i][5][7]),
        .io_output_5_8(mems_output[i][5][8]),
        .io_output_5_9(mems_output[i][5][9]),
        .io_output_5_10(mems_output[i][5][10]),
        .io_output_5_11(mems_output[i][5][11]),
        .io_output_5_12(mems_output[i][5][12]),
        .io_output_5_13(mems_output[i][5][13]),
        .io_output_5_14(mems_output[i][5][14]),
        .io_output_5_15(mems_output[i][5][15]),
        .io_output_5_16(mems_output[i][5][16]),
        .io_output_5_17(mems_output[i][5][17]),
        .io_output_5_18(mems_output[i][5][18]),
        .io_output_5_19(mems_output[i][5][19]),
        .io_output_5_20(mems_output[i][5][20]),
        .io_output_5_21(mems_output[i][5][21]),
        .io_output_5_22(mems_output[i][5][22]),
        .io_output_5_23(mems_output[i][5][23]),
        .io_output_5_24(mems_output[i][5][24]),
        .io_output_5_25(mems_output[i][5][25]),
        .io_output_5_26(mems_output[i][5][26]),
        .io_output_5_27(mems_output[i][5][27]),
        .io_output_5_28(mems_output[i][5][28]),
        .io_output_5_29(mems_output[i][5][29]),
        .io_output_5_30(mems_output[i][5][30]),
        .io_output_5_31(mems_output[i][5][31]),
        .io_output_6_0(mems_output[i][6][0]),
        .io_output_6_1(mems_output[i][6][1]),
        .io_output_6_2(mems_output[i][6][2]),
        .io_output_6_3(mems_output[i][6][3]),
        .io_output_6_4(mems_output[i][6][4]),
        .io_output_6_5(mems_output[i][6][5]),
        .io_output_6_6(mems_output[i][6][6]),
        .io_output_6_7(mems_output[i][6][7]),
        .io_output_6_8(mems_output[i][6][8]),
        .io_output_6_9(mems_output[i][6][9]),
        .io_output_6_10(mems_output[i][6][10]),
        .io_output_6_11(mems_output[i][6][11]),
        .io_output_6_12(mems_output[i][6][12]),
        .io_output_6_13(mems_output[i][6][13]),
        .io_output_6_14(mems_output[i][6][14]),
        .io_output_6_15(mems_output[i][6][15]),
        .io_output_6_16(mems_output[i][6][16]),
        .io_output_6_17(mems_output[i][6][17]),
        .io_output_6_18(mems_output[i][6][18]),
        .io_output_6_19(mems_output[i][6][19]),
        .io_output_6_20(mems_output[i][6][20]),
        .io_output_6_21(mems_output[i][6][21]),
        .io_output_6_22(mems_output[i][6][22]),
        .io_output_6_23(mems_output[i][6][23]),
        .io_output_6_24(mems_output[i][6][24]),
        .io_output_6_25(mems_output[i][6][25]),
        .io_output_6_26(mems_output[i][6][26]),
        .io_output_6_27(mems_output[i][6][27]),
        .io_output_6_28(mems_output[i][6][28]),
        .io_output_6_29(mems_output[i][6][29]),
        .io_output_6_30(mems_output[i][6][30]),
        .io_output_6_31(mems_output[i][6][31]),
        .io_output_7_0(mems_output[i][7][0]),
        .io_output_7_1(mems_output[i][7][1]),
        .io_output_7_2(mems_output[i][7][2]),
        .io_output_7_3(mems_output[i][7][3]),
        .io_output_7_4(mems_output[i][7][4]),
        .io_output_7_5(mems_output[i][7][5]),
        .io_output_7_6(mems_output[i][7][6]),
        .io_output_7_7(mems_output[i][7][7]),
        .io_output_7_8(mems_output[i][7][8]),
        .io_output_7_9(mems_output[i][7][9]),
        .io_output_7_10(mems_output[i][7][10]),
        .io_output_7_11(mems_output[i][7][11]),
        .io_output_7_12(mems_output[i][7][12]),
        .io_output_7_13(mems_output[i][7][13]),
        .io_output_7_14(mems_output[i][7][14]),
        .io_output_7_15(mems_output[i][7][15]),
        .io_output_7_16(mems_output[i][7][16]),
        .io_output_7_17(mems_output[i][7][17]),
        .io_output_7_18(mems_output[i][7][18]),
        .io_output_7_19(mems_output[i][7][19]),
        .io_output_7_20(mems_output[i][7][20]),
        .io_output_7_21(mems_output[i][7][21]),
        .io_output_7_22(mems_output[i][7][22]),
        .io_output_7_23(mems_output[i][7][23]),
        .io_output_7_24(mems_output[i][7][24]),
        .io_output_7_25(mems_output[i][7][25]),
        .io_output_7_26(mems_output[i][7][26]),
        .io_output_7_27(mems_output[i][7][27]),
        .io_output_7_28(mems_output[i][7][28]),
        .io_output_7_29(mems_output[i][7][29]),
        .io_output_7_30(mems_output[i][7][30]),
        .io_output_7_31(mems_output[i][7][31]),
        .io_output_8_0(mems_output[i][8][0]),
        .io_output_8_1(mems_output[i][8][1]),
        .io_output_8_2(mems_output[i][8][2]),
        .io_output_8_3(mems_output[i][8][3]),
        .io_output_8_4(mems_output[i][8][4]),
        .io_output_8_5(mems_output[i][8][5]),
        .io_output_8_6(mems_output[i][8][6]),
        .io_output_8_7(mems_output[i][8][7]),
        .io_output_8_8(mems_output[i][8][8]),
        .io_output_8_9(mems_output[i][8][9]),
        .io_output_8_10(mems_output[i][8][10]),
        .io_output_8_11(mems_output[i][8][11]),
        .io_output_8_12(mems_output[i][8][12]),
        .io_output_8_13(mems_output[i][8][13]),
        .io_output_8_14(mems_output[i][8][14]),
        .io_output_8_15(mems_output[i][8][15]),
        .io_output_8_16(mems_output[i][8][16]),
        .io_output_8_17(mems_output[i][8][17]),
        .io_output_8_18(mems_output[i][8][18]),
        .io_output_8_19(mems_output[i][8][19]),
        .io_output_8_20(mems_output[i][8][20]),
        .io_output_8_21(mems_output[i][8][21]),
        .io_output_8_22(mems_output[i][8][22]),
        .io_output_8_23(mems_output[i][8][23]),
        .io_output_8_24(mems_output[i][8][24]),
        .io_output_8_25(mems_output[i][8][25]),
        .io_output_8_26(mems_output[i][8][26]),
        .io_output_8_27(mems_output[i][8][27]),
        .io_output_8_28(mems_output[i][8][28]),
        .io_output_8_29(mems_output[i][8][29]),
        .io_output_8_30(mems_output[i][8][30]),
        .io_output_8_31(mems_output[i][8][31]),
        .io_output_9_0(mems_output[i][9][0]),
        .io_output_9_1(mems_output[i][9][1]),
        .io_output_9_2(mems_output[i][9][2]),
        .io_output_9_3(mems_output[i][9][3]),
        .io_output_9_4(mems_output[i][9][4]),
        .io_output_9_5(mems_output[i][9][5]),
        .io_output_9_6(mems_output[i][9][6]),
        .io_output_9_7(mems_output[i][9][7]),
        .io_output_9_8(mems_output[i][9][8]),
        .io_output_9_9(mems_output[i][9][9]),
        .io_output_9_10(mems_output[i][9][10]),
        .io_output_9_11(mems_output[i][9][11]),
        .io_output_9_12(mems_output[i][9][12]),
        .io_output_9_13(mems_output[i][9][13]),
        .io_output_9_14(mems_output[i][9][14]),
        .io_output_9_15(mems_output[i][9][15]),
        .io_output_9_16(mems_output[i][9][16]),
        .io_output_9_17(mems_output[i][9][17]),
        .io_output_9_18(mems_output[i][9][18]),
        .io_output_9_19(mems_output[i][9][19]),
        .io_output_9_20(mems_output[i][9][20]),
        .io_output_9_21(mems_output[i][9][21]),
        .io_output_9_22(mems_output[i][9][22]),
        .io_output_9_23(mems_output[i][9][23]),
        .io_output_9_24(mems_output[i][9][24]),
        .io_output_9_25(mems_output[i][9][25]),
        .io_output_9_26(mems_output[i][9][26]),
        .io_output_9_27(mems_output[i][9][27]),
        .io_output_9_28(mems_output[i][9][28]),
        .io_output_9_29(mems_output[i][9][29]),
        .io_output_9_30(mems_output[i][9][30]),
        .io_output_9_31(mems_output[i][9][31]),
        .io_output_10_0(mems_output[i][10][0]),
        .io_output_10_1(mems_output[i][10][1]),
        .io_output_10_2(mems_output[i][10][2]),
        .io_output_10_3(mems_output[i][10][3]),
        .io_output_10_4(mems_output[i][10][4]),
        .io_output_10_5(mems_output[i][10][5]),
        .io_output_10_6(mems_output[i][10][6]),
        .io_output_10_7(mems_output[i][10][7]),
        .io_output_10_8(mems_output[i][10][8]),
        .io_output_10_9(mems_output[i][10][9]),
        .io_output_10_10(mems_output[i][10][10]),
        .io_output_10_11(mems_output[i][10][11]),
        .io_output_10_12(mems_output[i][10][12]),
        .io_output_10_13(mems_output[i][10][13]),
        .io_output_10_14(mems_output[i][10][14]),
        .io_output_10_15(mems_output[i][10][15]),
        .io_output_10_16(mems_output[i][10][16]),
        .io_output_10_17(mems_output[i][10][17]),
        .io_output_10_18(mems_output[i][10][18]),
        .io_output_10_19(mems_output[i][10][19]),
        .io_output_10_20(mems_output[i][10][20]),
        .io_output_10_21(mems_output[i][10][21]),
        .io_output_10_22(mems_output[i][10][22]),
        .io_output_10_23(mems_output[i][10][23]),
        .io_output_10_24(mems_output[i][10][24]),
        .io_output_10_25(mems_output[i][10][25]),
        .io_output_10_26(mems_output[i][10][26]),
        .io_output_10_27(mems_output[i][10][27]),
        .io_output_10_28(mems_output[i][10][28]),
        .io_output_10_29(mems_output[i][10][29]),
        .io_output_10_30(mems_output[i][10][30]),
        .io_output_10_31(mems_output[i][10][31]),
        .io_output_11_0(mems_output[i][11][0]),
        .io_output_11_1(mems_output[i][11][1]),
        .io_output_11_2(mems_output[i][11][2]),
        .io_output_11_3(mems_output[i][11][3]),
        .io_output_11_4(mems_output[i][11][4]),
        .io_output_11_5(mems_output[i][11][5]),
        .io_output_11_6(mems_output[i][11][6]),
        .io_output_11_7(mems_output[i][11][7]),
        .io_output_11_8(mems_output[i][11][8]),
        .io_output_11_9(mems_output[i][11][9]),
        .io_output_11_10(mems_output[i][11][10]),
        .io_output_11_11(mems_output[i][11][11]),
        .io_output_11_12(mems_output[i][11][12]),
        .io_output_11_13(mems_output[i][11][13]),
        .io_output_11_14(mems_output[i][11][14]),
        .io_output_11_15(mems_output[i][11][15]),
        .io_output_11_16(mems_output[i][11][16]),
        .io_output_11_17(mems_output[i][11][17]),
        .io_output_11_18(mems_output[i][11][18]),
        .io_output_11_19(mems_output[i][11][19]),
        .io_output_11_20(mems_output[i][11][20]),
        .io_output_11_21(mems_output[i][11][21]),
        .io_output_11_22(mems_output[i][11][22]),
        .io_output_11_23(mems_output[i][11][23]),
        .io_output_11_24(mems_output[i][11][24]),
        .io_output_11_25(mems_output[i][11][25]),
        .io_output_11_26(mems_output[i][11][26]),
        .io_output_11_27(mems_output[i][11][27]),
        .io_output_11_28(mems_output[i][11][28]),
        .io_output_11_29(mems_output[i][11][29]),
        .io_output_11_30(mems_output[i][11][30]),
        .io_output_11_31(mems_output[i][11][31]),
        .io_output_12_0(mems_output[i][12][0]),
        .io_output_12_1(mems_output[i][12][1]),
        .io_output_12_2(mems_output[i][12][2]),
        .io_output_12_3(mems_output[i][12][3]),
        .io_output_12_4(mems_output[i][12][4]),
        .io_output_12_5(mems_output[i][12][5]),
        .io_output_12_6(mems_output[i][12][6]),
        .io_output_12_7(mems_output[i][12][7]),
        .io_output_12_8(mems_output[i][12][8]),
        .io_output_12_9(mems_output[i][12][9]),
        .io_output_12_10(mems_output[i][12][10]),
        .io_output_12_11(mems_output[i][12][11]),
        .io_output_12_12(mems_output[i][12][12]),
        .io_output_12_13(mems_output[i][12][13]),
        .io_output_12_14(mems_output[i][12][14]),
        .io_output_12_15(mems_output[i][12][15]),
        .io_output_12_16(mems_output[i][12][16]),
        .io_output_12_17(mems_output[i][12][17]),
        .io_output_12_18(mems_output[i][12][18]),
        .io_output_12_19(mems_output[i][12][19]),
        .io_output_12_20(mems_output[i][12][20]),
        .io_output_12_21(mems_output[i][12][21]),
        .io_output_12_22(mems_output[i][12][22]),
        .io_output_12_23(mems_output[i][12][23]),
        .io_output_12_24(mems_output[i][12][24]),
        .io_output_12_25(mems_output[i][12][25]),
        .io_output_12_26(mems_output[i][12][26]),
        .io_output_12_27(mems_output[i][12][27]),
        .io_output_12_28(mems_output[i][12][28]),
        .io_output_12_29(mems_output[i][12][29]),
        .io_output_12_30(mems_output[i][12][30]),
        .io_output_12_31(mems_output[i][12][31]),
        .io_output_13_0(mems_output[i][13][0]),
        .io_output_13_1(mems_output[i][13][1]),
        .io_output_13_2(mems_output[i][13][2]),
        .io_output_13_3(mems_output[i][13][3]),
        .io_output_13_4(mems_output[i][13][4]),
        .io_output_13_5(mems_output[i][13][5]),
        .io_output_13_6(mems_output[i][13][6]),
        .io_output_13_7(mems_output[i][13][7]),
        .io_output_13_8(mems_output[i][13][8]),
        .io_output_13_9(mems_output[i][13][9]),
        .io_output_13_10(mems_output[i][13][10]),
        .io_output_13_11(mems_output[i][13][11]),
        .io_output_13_12(mems_output[i][13][12]),
        .io_output_13_13(mems_output[i][13][13]),
        .io_output_13_14(mems_output[i][13][14]),
        .io_output_13_15(mems_output[i][13][15]),
        .io_output_13_16(mems_output[i][13][16]),
        .io_output_13_17(mems_output[i][13][17]),
        .io_output_13_18(mems_output[i][13][18]),
        .io_output_13_19(mems_output[i][13][19]),
        .io_output_13_20(mems_output[i][13][20]),
        .io_output_13_21(mems_output[i][13][21]),
        .io_output_13_22(mems_output[i][13][22]),
        .io_output_13_23(mems_output[i][13][23]),
        .io_output_13_24(mems_output[i][13][24]),
        .io_output_13_25(mems_output[i][13][25]),
        .io_output_13_26(mems_output[i][13][26]),
        .io_output_13_27(mems_output[i][13][27]),
        .io_output_13_28(mems_output[i][13][28]),
        .io_output_13_29(mems_output[i][13][29]),
        .io_output_13_30(mems_output[i][13][30]),
        .io_output_13_31(mems_output[i][13][31]),
        .io_output_14_0(mems_output[i][14][0]),
        .io_output_14_1(mems_output[i][14][1]),
        .io_output_14_2(mems_output[i][14][2]),
        .io_output_14_3(mems_output[i][14][3]),
        .io_output_14_4(mems_output[i][14][4]),
        .io_output_14_5(mems_output[i][14][5]),
        .io_output_14_6(mems_output[i][14][6]),
        .io_output_14_7(mems_output[i][14][7]),
        .io_output_14_8(mems_output[i][14][8]),
        .io_output_14_9(mems_output[i][14][9]),
        .io_output_14_10(mems_output[i][14][10]),
        .io_output_14_11(mems_output[i][14][11]),
        .io_output_14_12(mems_output[i][14][12]),
        .io_output_14_13(mems_output[i][14][13]),
        .io_output_14_14(mems_output[i][14][14]),
        .io_output_14_15(mems_output[i][14][15]),
        .io_output_14_16(mems_output[i][14][16]),
        .io_output_14_17(mems_output[i][14][17]),
        .io_output_14_18(mems_output[i][14][18]),
        .io_output_14_19(mems_output[i][14][19]),
        .io_output_14_20(mems_output[i][14][20]),
        .io_output_14_21(mems_output[i][14][21]),
        .io_output_14_22(mems_output[i][14][22]),
        .io_output_14_23(mems_output[i][14][23]),
        .io_output_14_24(mems_output[i][14][24]),
        .io_output_14_25(mems_output[i][14][25]),
        .io_output_14_26(mems_output[i][14][26]),
        .io_output_14_27(mems_output[i][14][27]),
        .io_output_14_28(mems_output[i][14][28]),
        .io_output_14_29(mems_output[i][14][29]),
        .io_output_14_30(mems_output[i][14][30]),
        .io_output_14_31(mems_output[i][14][31]),
        .io_output_15_0(mems_output[i][15][0]),
        .io_output_15_1(mems_output[i][15][1]),
        .io_output_15_2(mems_output[i][15][2]),
        .io_output_15_3(mems_output[i][15][3]),
        .io_output_15_4(mems_output[i][15][4]),
        .io_output_15_5(mems_output[i][15][5]),
        .io_output_15_6(mems_output[i][15][6]),
        .io_output_15_7(mems_output[i][15][7]),
        .io_output_15_8(mems_output[i][15][8]),
        .io_output_15_9(mems_output[i][15][9]),
        .io_output_15_10(mems_output[i][15][10]),
        .io_output_15_11(mems_output[i][15][11]),
        .io_output_15_12(mems_output[i][15][12]),
        .io_output_15_13(mems_output[i][15][13]),
        .io_output_15_14(mems_output[i][15][14]),
        .io_output_15_15(mems_output[i][15][15]),
        .io_output_15_16(mems_output[i][15][16]),
        .io_output_15_17(mems_output[i][15][17]),
        .io_output_15_18(mems_output[i][15][18]),
        .io_output_15_19(mems_output[i][15][19]),
        .io_output_15_20(mems_output[i][15][20]),
        .io_output_15_21(mems_output[i][15][21]),
        .io_output_15_22(mems_output[i][15][22]),
        .io_output_15_23(mems_output[i][15][23]),
        .io_output_15_24(mems_output[i][15][24]),
        .io_output_15_25(mems_output[i][15][25]),
        .io_output_15_26(mems_output[i][15][26]),
        .io_output_15_27(mems_output[i][15][27]),
        .io_output_15_28(mems_output[i][15][28]),
        .io_output_15_29(mems_output[i][15][29]),
        .io_output_15_30(mems_output[i][15][30]),
        .io_output_15_31(mems_output[i][15][31]),
        .io_output_16_0(mems_output[i][16][0]),
        .io_output_16_1(mems_output[i][16][1]),
        .io_output_16_2(mems_output[i][16][2]),
        .io_output_16_3(mems_output[i][16][3]),
        .io_output_16_4(mems_output[i][16][4]),
        .io_output_16_5(mems_output[i][16][5]),
        .io_output_16_6(mems_output[i][16][6]),
        .io_output_16_7(mems_output[i][16][7]),
        .io_output_16_8(mems_output[i][16][8]),
        .io_output_16_9(mems_output[i][16][9]),
        .io_output_16_10(mems_output[i][16][10]),
        .io_output_16_11(mems_output[i][16][11]),
        .io_output_16_12(mems_output[i][16][12]),
        .io_output_16_13(mems_output[i][16][13]),
        .io_output_16_14(mems_output[i][16][14]),
        .io_output_16_15(mems_output[i][16][15]),
        .io_output_16_16(mems_output[i][16][16]),
        .io_output_16_17(mems_output[i][16][17]),
        .io_output_16_18(mems_output[i][16][18]),
        .io_output_16_19(mems_output[i][16][19]),
        .io_output_16_20(mems_output[i][16][20]),
        .io_output_16_21(mems_output[i][16][21]),
        .io_output_16_22(mems_output[i][16][22]),
        .io_output_16_23(mems_output[i][16][23]),
        .io_output_16_24(mems_output[i][16][24]),
        .io_output_16_25(mems_output[i][16][25]),
        .io_output_16_26(mems_output[i][16][26]),
        .io_output_16_27(mems_output[i][16][27]),
        .io_output_16_28(mems_output[i][16][28]),
        .io_output_16_29(mems_output[i][16][29]),
        .io_output_16_30(mems_output[i][16][30]),
        .io_output_16_31(mems_output[i][16][31]),
        .io_output_17_0(mems_output[i][17][0]),
        .io_output_17_1(mems_output[i][17][1]),
        .io_output_17_2(mems_output[i][17][2]),
        .io_output_17_3(mems_output[i][17][3]),
        .io_output_17_4(mems_output[i][17][4]),
        .io_output_17_5(mems_output[i][17][5]),
        .io_output_17_6(mems_output[i][17][6]),
        .io_output_17_7(mems_output[i][17][7]),
        .io_output_17_8(mems_output[i][17][8]),
        .io_output_17_9(mems_output[i][17][9]),
        .io_output_17_10(mems_output[i][17][10]),
        .io_output_17_11(mems_output[i][17][11]),
        .io_output_17_12(mems_output[i][17][12]),
        .io_output_17_13(mems_output[i][17][13]),
        .io_output_17_14(mems_output[i][17][14]),
        .io_output_17_15(mems_output[i][17][15]),
        .io_output_17_16(mems_output[i][17][16]),
        .io_output_17_17(mems_output[i][17][17]),
        .io_output_17_18(mems_output[i][17][18]),
        .io_output_17_19(mems_output[i][17][19]),
        .io_output_17_20(mems_output[i][17][20]),
        .io_output_17_21(mems_output[i][17][21]),
        .io_output_17_22(mems_output[i][17][22]),
        .io_output_17_23(mems_output[i][17][23]),
        .io_output_17_24(mems_output[i][17][24]),
        .io_output_17_25(mems_output[i][17][25]),
        .io_output_17_26(mems_output[i][17][26]),
        .io_output_17_27(mems_output[i][17][27]),
        .io_output_17_28(mems_output[i][17][28]),
        .io_output_17_29(mems_output[i][17][29]),
        .io_output_17_30(mems_output[i][17][30]),
        .io_output_17_31(mems_output[i][17][31]),
        .io_output_18_0(mems_output[i][18][0]),
        .io_output_18_1(mems_output[i][18][1]),
        .io_output_18_2(mems_output[i][18][2]),
        .io_output_18_3(mems_output[i][18][3]),
        .io_output_18_4(mems_output[i][18][4]),
        .io_output_18_5(mems_output[i][18][5]),
        .io_output_18_6(mems_output[i][18][6]),
        .io_output_18_7(mems_output[i][18][7]),
        .io_output_18_8(mems_output[i][18][8]),
        .io_output_18_9(mems_output[i][18][9]),
        .io_output_18_10(mems_output[i][18][10]),
        .io_output_18_11(mems_output[i][18][11]),
        .io_output_18_12(mems_output[i][18][12]),
        .io_output_18_13(mems_output[i][18][13]),
        .io_output_18_14(mems_output[i][18][14]),
        .io_output_18_15(mems_output[i][18][15]),
        .io_output_18_16(mems_output[i][18][16]),
        .io_output_18_17(mems_output[i][18][17]),
        .io_output_18_18(mems_output[i][18][18]),
        .io_output_18_19(mems_output[i][18][19]),
        .io_output_18_20(mems_output[i][18][20]),
        .io_output_18_21(mems_output[i][18][21]),
        .io_output_18_22(mems_output[i][18][22]),
        .io_output_18_23(mems_output[i][18][23]),
        .io_output_18_24(mems_output[i][18][24]),
        .io_output_18_25(mems_output[i][18][25]),
        .io_output_18_26(mems_output[i][18][26]),
        .io_output_18_27(mems_output[i][18][27]),
        .io_output_18_28(mems_output[i][18][28]),
        .io_output_18_29(mems_output[i][18][29]),
        .io_output_18_30(mems_output[i][18][30]),
        .io_output_18_31(mems_output[i][18][31]),
        .io_output_19_0(mems_output[i][19][0]),
        .io_output_19_1(mems_output[i][19][1]),
        .io_output_19_2(mems_output[i][19][2]),
        .io_output_19_3(mems_output[i][19][3]),
        .io_output_19_4(mems_output[i][19][4]),
        .io_output_19_5(mems_output[i][19][5]),
        .io_output_19_6(mems_output[i][19][6]),
        .io_output_19_7(mems_output[i][19][7]),
        .io_output_19_8(mems_output[i][19][8]),
        .io_output_19_9(mems_output[i][19][9]),
        .io_output_19_10(mems_output[i][19][10]),
        .io_output_19_11(mems_output[i][19][11]),
        .io_output_19_12(mems_output[i][19][12]),
        .io_output_19_13(mems_output[i][19][13]),
        .io_output_19_14(mems_output[i][19][14]),
        .io_output_19_15(mems_output[i][19][15]),
        .io_output_19_16(mems_output[i][19][16]),
        .io_output_19_17(mems_output[i][19][17]),
        .io_output_19_18(mems_output[i][19][18]),
        .io_output_19_19(mems_output[i][19][19]),
        .io_output_19_20(mems_output[i][19][20]),
        .io_output_19_21(mems_output[i][19][21]),
        .io_output_19_22(mems_output[i][19][22]),
        .io_output_19_23(mems_output[i][19][23]),
        .io_output_19_24(mems_output[i][19][24]),
        .io_output_19_25(mems_output[i][19][25]),
        .io_output_19_26(mems_output[i][19][26]),
        .io_output_19_27(mems_output[i][19][27]),
        .io_output_19_28(mems_output[i][19][28]),
        .io_output_19_29(mems_output[i][19][29]),
        .io_output_19_30(mems_output[i][19][30]),
        .io_output_19_31(mems_output[i][19][31]),
        .io_output_20_0(mems_output[i][20][0]),
        .io_output_20_1(mems_output[i][20][1]),
        .io_output_20_2(mems_output[i][20][2]),
        .io_output_20_3(mems_output[i][20][3]),
        .io_output_20_4(mems_output[i][20][4]),
        .io_output_20_5(mems_output[i][20][5]),
        .io_output_20_6(mems_output[i][20][6]),
        .io_output_20_7(mems_output[i][20][7]),
        .io_output_20_8(mems_output[i][20][8]),
        .io_output_20_9(mems_output[i][20][9]),
        .io_output_20_10(mems_output[i][20][10]),
        .io_output_20_11(mems_output[i][20][11]),
        .io_output_20_12(mems_output[i][20][12]),
        .io_output_20_13(mems_output[i][20][13]),
        .io_output_20_14(mems_output[i][20][14]),
        .io_output_20_15(mems_output[i][20][15]),
        .io_output_20_16(mems_output[i][20][16]),
        .io_output_20_17(mems_output[i][20][17]),
        .io_output_20_18(mems_output[i][20][18]),
        .io_output_20_19(mems_output[i][20][19]),
        .io_output_20_20(mems_output[i][20][20]),
        .io_output_20_21(mems_output[i][20][21]),
        .io_output_20_22(mems_output[i][20][22]),
        .io_output_20_23(mems_output[i][20][23]),
        .io_output_20_24(mems_output[i][20][24]),
        .io_output_20_25(mems_output[i][20][25]),
        .io_output_20_26(mems_output[i][20][26]),
        .io_output_20_27(mems_output[i][20][27]),
        .io_output_20_28(mems_output[i][20][28]),
        .io_output_20_29(mems_output[i][20][29]),
        .io_output_20_30(mems_output[i][20][30]),
        .io_output_20_31(mems_output[i][20][31]),
        .io_output_21_0(mems_output[i][21][0]),
        .io_output_21_1(mems_output[i][21][1]),
        .io_output_21_2(mems_output[i][21][2]),
        .io_output_21_3(mems_output[i][21][3]),
        .io_output_21_4(mems_output[i][21][4]),
        .io_output_21_5(mems_output[i][21][5]),
        .io_output_21_6(mems_output[i][21][6]),
        .io_output_21_7(mems_output[i][21][7]),
        .io_output_21_8(mems_output[i][21][8]),
        .io_output_21_9(mems_output[i][21][9]),
        .io_output_21_10(mems_output[i][21][10]),
        .io_output_21_11(mems_output[i][21][11]),
        .io_output_21_12(mems_output[i][21][12]),
        .io_output_21_13(mems_output[i][21][13]),
        .io_output_21_14(mems_output[i][21][14]),
        .io_output_21_15(mems_output[i][21][15]),
        .io_output_21_16(mems_output[i][21][16]),
        .io_output_21_17(mems_output[i][21][17]),
        .io_output_21_18(mems_output[i][21][18]),
        .io_output_21_19(mems_output[i][21][19]),
        .io_output_21_20(mems_output[i][21][20]),
        .io_output_21_21(mems_output[i][21][21]),
        .io_output_21_22(mems_output[i][21][22]),
        .io_output_21_23(mems_output[i][21][23]),
        .io_output_21_24(mems_output[i][21][24]),
        .io_output_21_25(mems_output[i][21][25]),
        .io_output_21_26(mems_output[i][21][26]),
        .io_output_21_27(mems_output[i][21][27]),
        .io_output_21_28(mems_output[i][21][28]),
        .io_output_21_29(mems_output[i][21][29]),
        .io_output_21_30(mems_output[i][21][30]),
        .io_output_21_31(mems_output[i][21][31]),
        .io_output_22_0(mems_output[i][22][0]),
        .io_output_22_1(mems_output[i][22][1]),
        .io_output_22_2(mems_output[i][22][2]),
        .io_output_22_3(mems_output[i][22][3]),
        .io_output_22_4(mems_output[i][22][4]),
        .io_output_22_5(mems_output[i][22][5]),
        .io_output_22_6(mems_output[i][22][6]),
        .io_output_22_7(mems_output[i][22][7]),
        .io_output_22_8(mems_output[i][22][8]),
        .io_output_22_9(mems_output[i][22][9]),
        .io_output_22_10(mems_output[i][22][10]),
        .io_output_22_11(mems_output[i][22][11]),
        .io_output_22_12(mems_output[i][22][12]),
        .io_output_22_13(mems_output[i][22][13]),
        .io_output_22_14(mems_output[i][22][14]),
        .io_output_22_15(mems_output[i][22][15]),
        .io_output_22_16(mems_output[i][22][16]),
        .io_output_22_17(mems_output[i][22][17]),
        .io_output_22_18(mems_output[i][22][18]),
        .io_output_22_19(mems_output[i][22][19]),
        .io_output_22_20(mems_output[i][22][20]),
        .io_output_22_21(mems_output[i][22][21]),
        .io_output_22_22(mems_output[i][22][22]),
        .io_output_22_23(mems_output[i][22][23]),
        .io_output_22_24(mems_output[i][22][24]),
        .io_output_22_25(mems_output[i][22][25]),
        .io_output_22_26(mems_output[i][22][26]),
        .io_output_22_27(mems_output[i][22][27]),
        .io_output_22_28(mems_output[i][22][28]),
        .io_output_22_29(mems_output[i][22][29]),
        .io_output_22_30(mems_output[i][22][30]),
        .io_output_22_31(mems_output[i][22][31]),
        .io_output_23_0(mems_output[i][23][0]),
        .io_output_23_1(mems_output[i][23][1]),
        .io_output_23_2(mems_output[i][23][2]),
        .io_output_23_3(mems_output[i][23][3]),
        .io_output_23_4(mems_output[i][23][4]),
        .io_output_23_5(mems_output[i][23][5]),
        .io_output_23_6(mems_output[i][23][6]),
        .io_output_23_7(mems_output[i][23][7]),
        .io_output_23_8(mems_output[i][23][8]),
        .io_output_23_9(mems_output[i][23][9]),
        .io_output_23_10(mems_output[i][23][10]),
        .io_output_23_11(mems_output[i][23][11]),
        .io_output_23_12(mems_output[i][23][12]),
        .io_output_23_13(mems_output[i][23][13]),
        .io_output_23_14(mems_output[i][23][14]),
        .io_output_23_15(mems_output[i][23][15]),
        .io_output_23_16(mems_output[i][23][16]),
        .io_output_23_17(mems_output[i][23][17]),
        .io_output_23_18(mems_output[i][23][18]),
        .io_output_23_19(mems_output[i][23][19]),
        .io_output_23_20(mems_output[i][23][20]),
        .io_output_23_21(mems_output[i][23][21]),
        .io_output_23_22(mems_output[i][23][22]),
        .io_output_23_23(mems_output[i][23][23]),
        .io_output_23_24(mems_output[i][23][24]),
        .io_output_23_25(mems_output[i][23][25]),
        .io_output_23_26(mems_output[i][23][26]),
        .io_output_23_27(mems_output[i][23][27]),
        .io_output_23_28(mems_output[i][23][28]),
        .io_output_23_29(mems_output[i][23][29]),
        .io_output_23_30(mems_output[i][23][30]),
        .io_output_23_31(mems_output[i][23][31]),
        .io_output_24_0(mems_output[i][24][0]),
        .io_output_24_1(mems_output[i][24][1]),
        .io_output_24_2(mems_output[i][24][2]),
        .io_output_24_3(mems_output[i][24][3]),
        .io_output_24_4(mems_output[i][24][4]),
        .io_output_24_5(mems_output[i][24][5]),
        .io_output_24_6(mems_output[i][24][6]),
        .io_output_24_7(mems_output[i][24][7]),
        .io_output_24_8(mems_output[i][24][8]),
        .io_output_24_9(mems_output[i][24][9]),
        .io_output_24_10(mems_output[i][24][10]),
        .io_output_24_11(mems_output[i][24][11]),
        .io_output_24_12(mems_output[i][24][12]),
        .io_output_24_13(mems_output[i][24][13]),
        .io_output_24_14(mems_output[i][24][14]),
        .io_output_24_15(mems_output[i][24][15]),
        .io_output_24_16(mems_output[i][24][16]),
        .io_output_24_17(mems_output[i][24][17]),
        .io_output_24_18(mems_output[i][24][18]),
        .io_output_24_19(mems_output[i][24][19]),
        .io_output_24_20(mems_output[i][24][20]),
        .io_output_24_21(mems_output[i][24][21]),
        .io_output_24_22(mems_output[i][24][22]),
        .io_output_24_23(mems_output[i][24][23]),
        .io_output_24_24(mems_output[i][24][24]),
        .io_output_24_25(mems_output[i][24][25]),
        .io_output_24_26(mems_output[i][24][26]),
        .io_output_24_27(mems_output[i][24][27]),
        .io_output_24_28(mems_output[i][24][28]),
        .io_output_24_29(mems_output[i][24][29]),
        .io_output_24_30(mems_output[i][24][30]),
        .io_output_24_31(mems_output[i][24][31]),
        .io_output_25_0(mems_output[i][25][0]),
        .io_output_25_1(mems_output[i][25][1]),
        .io_output_25_2(mems_output[i][25][2]),
        .io_output_25_3(mems_output[i][25][3]),
        .io_output_25_4(mems_output[i][25][4]),
        .io_output_25_5(mems_output[i][25][5]),
        .io_output_25_6(mems_output[i][25][6]),
        .io_output_25_7(mems_output[i][25][7]),
        .io_output_25_8(mems_output[i][25][8]),
        .io_output_25_9(mems_output[i][25][9]),
        .io_output_25_10(mems_output[i][25][10]),
        .io_output_25_11(mems_output[i][25][11]),
        .io_output_25_12(mems_output[i][25][12]),
        .io_output_25_13(mems_output[i][25][13]),
        .io_output_25_14(mems_output[i][25][14]),
        .io_output_25_15(mems_output[i][25][15]),
        .io_output_25_16(mems_output[i][25][16]),
        .io_output_25_17(mems_output[i][25][17]),
        .io_output_25_18(mems_output[i][25][18]),
        .io_output_25_19(mems_output[i][25][19]),
        .io_output_25_20(mems_output[i][25][20]),
        .io_output_25_21(mems_output[i][25][21]),
        .io_output_25_22(mems_output[i][25][22]),
        .io_output_25_23(mems_output[i][25][23]),
        .io_output_25_24(mems_output[i][25][24]),
        .io_output_25_25(mems_output[i][25][25]),
        .io_output_25_26(mems_output[i][25][26]),
        .io_output_25_27(mems_output[i][25][27]),
        .io_output_25_28(mems_output[i][25][28]),
        .io_output_25_29(mems_output[i][25][29]),
        .io_output_25_30(mems_output[i][25][30]),
        .io_output_25_31(mems_output[i][25][31]),
        .io_output_26_0(mems_output[i][26][0]),
        .io_output_26_1(mems_output[i][26][1]),
        .io_output_26_2(mems_output[i][26][2]),
        .io_output_26_3(mems_output[i][26][3]),
        .io_output_26_4(mems_output[i][26][4]),
        .io_output_26_5(mems_output[i][26][5]),
        .io_output_26_6(mems_output[i][26][6]),
        .io_output_26_7(mems_output[i][26][7]),
        .io_output_26_8(mems_output[i][26][8]),
        .io_output_26_9(mems_output[i][26][9]),
        .io_output_26_10(mems_output[i][26][10]),
        .io_output_26_11(mems_output[i][26][11]),
        .io_output_26_12(mems_output[i][26][12]),
        .io_output_26_13(mems_output[i][26][13]),
        .io_output_26_14(mems_output[i][26][14]),
        .io_output_26_15(mems_output[i][26][15]),
        .io_output_26_16(mems_output[i][26][16]),
        .io_output_26_17(mems_output[i][26][17]),
        .io_output_26_18(mems_output[i][26][18]),
        .io_output_26_19(mems_output[i][26][19]),
        .io_output_26_20(mems_output[i][26][20]),
        .io_output_26_21(mems_output[i][26][21]),
        .io_output_26_22(mems_output[i][26][22]),
        .io_output_26_23(mems_output[i][26][23]),
        .io_output_26_24(mems_output[i][26][24]),
        .io_output_26_25(mems_output[i][26][25]),
        .io_output_26_26(mems_output[i][26][26]),
        .io_output_26_27(mems_output[i][26][27]),
        .io_output_26_28(mems_output[i][26][28]),
        .io_output_26_29(mems_output[i][26][29]),
        .io_output_26_30(mems_output[i][26][30]),
        .io_output_26_31(mems_output[i][26][31]),
        .io_output_27_0(mems_output[i][27][0]),
        .io_output_27_1(mems_output[i][27][1]),
        .io_output_27_2(mems_output[i][27][2]),
        .io_output_27_3(mems_output[i][27][3]),
        .io_output_27_4(mems_output[i][27][4]),
        .io_output_27_5(mems_output[i][27][5]),
        .io_output_27_6(mems_output[i][27][6]),
        .io_output_27_7(mems_output[i][27][7]),
        .io_output_27_8(mems_output[i][27][8]),
        .io_output_27_9(mems_output[i][27][9]),
        .io_output_27_10(mems_output[i][27][10]),
        .io_output_27_11(mems_output[i][27][11]),
        .io_output_27_12(mems_output[i][27][12]),
        .io_output_27_13(mems_output[i][27][13]),
        .io_output_27_14(mems_output[i][27][14]),
        .io_output_27_15(mems_output[i][27][15]),
        .io_output_27_16(mems_output[i][27][16]),
        .io_output_27_17(mems_output[i][27][17]),
        .io_output_27_18(mems_output[i][27][18]),
        .io_output_27_19(mems_output[i][27][19]),
        .io_output_27_20(mems_output[i][27][20]),
        .io_output_27_21(mems_output[i][27][21]),
        .io_output_27_22(mems_output[i][27][22]),
        .io_output_27_23(mems_output[i][27][23]),
        .io_output_27_24(mems_output[i][27][24]),
        .io_output_27_25(mems_output[i][27][25]),
        .io_output_27_26(mems_output[i][27][26]),
        .io_output_27_27(mems_output[i][27][27]),
        .io_output_27_28(mems_output[i][27][28]),
        .io_output_27_29(mems_output[i][27][29]),
        .io_output_27_30(mems_output[i][27][30]),
        .io_output_27_31(mems_output[i][27][31]),
        .io_output_28_0(mems_output[i][28][0]),
        .io_output_28_1(mems_output[i][28][1]),
        .io_output_28_2(mems_output[i][28][2]),
        .io_output_28_3(mems_output[i][28][3]),
        .io_output_28_4(mems_output[i][28][4]),
        .io_output_28_5(mems_output[i][28][5]),
        .io_output_28_6(mems_output[i][28][6]),
        .io_output_28_7(mems_output[i][28][7]),
        .io_output_28_8(mems_output[i][28][8]),
        .io_output_28_9(mems_output[i][28][9]),
        .io_output_28_10(mems_output[i][28][10]),
        .io_output_28_11(mems_output[i][28][11]),
        .io_output_28_12(mems_output[i][28][12]),
        .io_output_28_13(mems_output[i][28][13]),
        .io_output_28_14(mems_output[i][28][14]),
        .io_output_28_15(mems_output[i][28][15]),
        .io_output_28_16(mems_output[i][28][16]),
        .io_output_28_17(mems_output[i][28][17]),
        .io_output_28_18(mems_output[i][28][18]),
        .io_output_28_19(mems_output[i][28][19]),
        .io_output_28_20(mems_output[i][28][20]),
        .io_output_28_21(mems_output[i][28][21]),
        .io_output_28_22(mems_output[i][28][22]),
        .io_output_28_23(mems_output[i][28][23]),
        .io_output_28_24(mems_output[i][28][24]),
        .io_output_28_25(mems_output[i][28][25]),
        .io_output_28_26(mems_output[i][28][26]),
        .io_output_28_27(mems_output[i][28][27]),
        .io_output_28_28(mems_output[i][28][28]),
        .io_output_28_29(mems_output[i][28][29]),
        .io_output_28_30(mems_output[i][28][30]),
        .io_output_28_31(mems_output[i][28][31]),
        .io_output_29_0(mems_output[i][29][0]),
        .io_output_29_1(mems_output[i][29][1]),
        .io_output_29_2(mems_output[i][29][2]),
        .io_output_29_3(mems_output[i][29][3]),
        .io_output_29_4(mems_output[i][29][4]),
        .io_output_29_5(mems_output[i][29][5]),
        .io_output_29_6(mems_output[i][29][6]),
        .io_output_29_7(mems_output[i][29][7]),
        .io_output_29_8(mems_output[i][29][8]),
        .io_output_29_9(mems_output[i][29][9]),
        .io_output_29_10(mems_output[i][29][10]),
        .io_output_29_11(mems_output[i][29][11]),
        .io_output_29_12(mems_output[i][29][12]),
        .io_output_29_13(mems_output[i][29][13]),
        .io_output_29_14(mems_output[i][29][14]),
        .io_output_29_15(mems_output[i][29][15]),
        .io_output_29_16(mems_output[i][29][16]),
        .io_output_29_17(mems_output[i][29][17]),
        .io_output_29_18(mems_output[i][29][18]),
        .io_output_29_19(mems_output[i][29][19]),
        .io_output_29_20(mems_output[i][29][20]),
        .io_output_29_21(mems_output[i][29][21]),
        .io_output_29_22(mems_output[i][29][22]),
        .io_output_29_23(mems_output[i][29][23]),
        .io_output_29_24(mems_output[i][29][24]),
        .io_output_29_25(mems_output[i][29][25]),
        .io_output_29_26(mems_output[i][29][26]),
        .io_output_29_27(mems_output[i][29][27]),
        .io_output_29_28(mems_output[i][29][28]),
        .io_output_29_29(mems_output[i][29][29]),
        .io_output_29_30(mems_output[i][29][30]),
        .io_output_29_31(mems_output[i][29][31]),
        .io_output_30_0(mems_output[i][30][0]),
        .io_output_30_1(mems_output[i][30][1]),
        .io_output_30_2(mems_output[i][30][2]),
        .io_output_30_3(mems_output[i][30][3]),
        .io_output_30_4(mems_output[i][30][4]),
        .io_output_30_5(mems_output[i][30][5]),
        .io_output_30_6(mems_output[i][30][6]),
        .io_output_30_7(mems_output[i][30][7]),
        .io_output_30_8(mems_output[i][30][8]),
        .io_output_30_9(mems_output[i][30][9]),
        .io_output_30_10(mems_output[i][30][10]),
        .io_output_30_11(mems_output[i][30][11]),
        .io_output_30_12(mems_output[i][30][12]),
        .io_output_30_13(mems_output[i][30][13]),
        .io_output_30_14(mems_output[i][30][14]),
        .io_output_30_15(mems_output[i][30][15]),
        .io_output_30_16(mems_output[i][30][16]),
        .io_output_30_17(mems_output[i][30][17]),
        .io_output_30_18(mems_output[i][30][18]),
        .io_output_30_19(mems_output[i][30][19]),
        .io_output_30_20(mems_output[i][30][20]),
        .io_output_30_21(mems_output[i][30][21]),
        .io_output_30_22(mems_output[i][30][22]),
        .io_output_30_23(mems_output[i][30][23]),
        .io_output_30_24(mems_output[i][30][24]),
        .io_output_30_25(mems_output[i][30][25]),
        .io_output_30_26(mems_output[i][30][26]),
        .io_output_30_27(mems_output[i][30][27]),
        .io_output_30_28(mems_output[i][30][28]),
        .io_output_30_29(mems_output[i][30][29]),
        .io_output_30_30(mems_output[i][30][30]),
        .io_output_30_31(mems_output[i][30][31]),
        .io_output_31_0(mems_output[i][31][0]),
        .io_output_31_1(mems_output[i][31][1]),
        .io_output_31_2(mems_output[i][31][2]),
        .io_output_31_3(mems_output[i][31][3]),
        .io_output_31_4(mems_output[i][31][4]),
        .io_output_31_5(mems_output[i][31][5]),
        .io_output_31_6(mems_output[i][31][6]),
        .io_output_31_7(mems_output[i][31][7]),
        .io_output_31_8(mems_output[i][31][8]),
        .io_output_31_9(mems_output[i][31][9]),
        .io_output_31_10(mems_output[i][31][10]),
        .io_output_31_11(mems_output[i][31][11]),
        .io_output_31_12(mems_output[i][31][12]),
        .io_output_31_13(mems_output[i][31][13]),
        .io_output_31_14(mems_output[i][31][14]),
        .io_output_31_15(mems_output[i][31][15]),
        .io_output_31_16(mems_output[i][31][16]),
        .io_output_31_17(mems_output[i][31][17]),
        .io_output_31_18(mems_output[i][31][18]),
        .io_output_31_19(mems_output[i][31][19]),
        .io_output_31_20(mems_output[i][31][20]),
        .io_output_31_21(mems_output[i][31][21]),
        .io_output_31_22(mems_output[i][31][22]),
        .io_output_31_23(mems_output[i][31][23]),
        .io_output_31_24(mems_output[i][31][24]),
        .io_output_31_25(mems_output[i][31][25]),
        .io_output_31_26(mems_output[i][31][26]),
        .io_output_31_27(mems_output[i][31][27]),
        .io_output_31_28(mems_output[i][31][28]),
        .io_output_31_29(mems_output[i][31][29]),
        .io_output_31_30(mems_output[i][31][30]),
        .io_output_31_31(mems_output[i][31][31])
    );
end endgenerate
//-----------------------------------------------------------------------------

//-----------------------------------------------------------------------------
// Include experiment file defined on command line 
//-----------------------------------------------------------------------------
`include `EXPERIMENT
//-----------------------------------------------------------------------------

//-----------------------------------------------------------------------------
// Execute test
//-----------------------------------------------------------------------------
//`ifdef CSVDATA
//int fd;
//always @(posedge bfm.i_clk) begin
//    if (bfm.o_decision_trigger) begin
//        bfm.dec_counter = bfm.dec_counter + 1;
//        $fdisplay(fd,"%d,%d,%d", bfm.dec_counter, bfm.o_heat_out, bfm.o_current_power);
//        //$display("Decision: %d", dec_counter);
//    end
//end
//`endif
    
initial begin
//`ifdef CSVDATA
//    // Open file for writing
//    fd = $fopen("data.csv", "w");
//    $fdisplay(fd, "decision,heat_code,power,ring_lambda");
//`endif

    // Pre experiment initialization
    // TODO

    run_experiment;

    $finish;

end
//-----------------------------------------------------------------------------

endmodule : top
